../../common/tb/prover_compute_w0_test.sv