../../common/rtl/verifier_compute_io.sv