../../common/rtl/verifier_layer.sv