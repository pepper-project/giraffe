../../common/tb/pergate_compute_gatefn_early_test.sv