../../common/rtl/verifier_compute_chi.sv