../../common/rtl/prover_shim_negate.sv