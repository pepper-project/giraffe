../../common/rtl/prover_compute_v_encollect.sv