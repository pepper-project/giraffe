../../common/tb/prover_interpolate_quadratic_test.sv