../../common/tb/prover_compute_v_late_gates_test.sv