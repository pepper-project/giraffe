../../common/rtl/prover_shuffle_early.sv