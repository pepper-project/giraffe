../../common/func/func_gateInNum.sv