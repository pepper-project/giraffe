../../common/tb/vpintf_test.sv