../../common/tb/verifier_compute_chi_dotp_test.sv