../../common/tb/prover_compute_chi_test.sv