../../common/rtl/prover_compute_chi.sv