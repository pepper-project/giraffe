../../common/tb/verifier_compute_beta_test.sv