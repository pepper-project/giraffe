../../common/tb/prover_compute_v_sr_test.sv