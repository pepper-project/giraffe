../../common/rtl/prover_compute_v_early_gatesbank.sv