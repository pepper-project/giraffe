../../common/tb/verifier_compute_chi_test.sv