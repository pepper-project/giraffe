../../common/rtl/prover_compute_h_accum.sv