../../common/rtl/prover_compute_v_srelem.sv