../../common/tb/prover_compute_v_encollect_test.sv