../../common/tb/verifier_compute_horner_test.sv