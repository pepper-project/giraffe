../../common/rtl/prover_compute_v_valsbank.sv