../../common/rtl/verifier_compute_chi_elem.sv