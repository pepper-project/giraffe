../../common/tb/lagrange_interpolate_test.sv