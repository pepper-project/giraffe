../../common/rtl/lagrange_coeffs.sv