../../common/tb/prover_compute_h_percopy_test.sv