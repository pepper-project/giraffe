../../common/tb/prover_lsb_posn_test.sv