../../common/rtl/prover_compute_h_parmux.sv