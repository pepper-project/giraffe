../../common/rtl/verifier_compute_chi_single.sv