../../common/rtl/verifier_compute_io_elem.sv