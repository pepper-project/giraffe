../../common/rtl/verifier_compute_wpreds.sv