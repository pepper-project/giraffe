../../common/rtl/prover_compute_v_late.sv