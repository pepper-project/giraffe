../../common/rtl/verifier_compute_io_elembank.sv