../../common/rtl/prover_compute_v_srbank.sv