../../common/rtl/verifier_compute_horner.sv