../../common/tb/verifier_layer_test.sv