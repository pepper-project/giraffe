../../common/rtl/pergate_compute_late.sv