../../common/rtl/prover_interpolate_cubic.sv