../../common/func/func_ithLagrangeCoeffs.sv