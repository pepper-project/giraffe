../../common/rtl/lagrange_interpolate.sv