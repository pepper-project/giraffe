../../common/tb/prover_shuffle_early_test.sv