../../common/rtl/prover_interpolate_qc.sv