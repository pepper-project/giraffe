../../common/rtl/computation_layer_elem.sv