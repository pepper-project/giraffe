../../common/tb/prover_compute_h_chi_test.sv