../../common/rtl/prover_interpolate_quadratic.sv