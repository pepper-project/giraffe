../../common/tb/prover_shim_test.sv