../../common/tb/verifier_adder_tree_test.sv