../../common/func/func_convertIntMtoL.sv