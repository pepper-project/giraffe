../../common/rtl/verifier_compute_beta.sv