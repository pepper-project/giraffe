../../common/tb/field_halve_test.sv