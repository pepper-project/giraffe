../../common/tb/verifier_compute_io_test.sv