../../common/func/func_leastSetBitPosn.sv