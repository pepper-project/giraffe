../../common/rtl/prover_compute_h_percopy.sv