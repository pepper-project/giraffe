../../common/rtl/field_halve.sv