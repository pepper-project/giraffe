../../common/tb/prover_compute_v_srbank_test.sv