../../common/rtl/pergate_compute_gatefn_early.sv