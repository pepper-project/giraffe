../../common/rtl/prover_compute_h_mulonly.sv