../../common/rtl/prover_compute_h_chi.sv