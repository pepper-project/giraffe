../../common/tb/verifier_compute_chi_single_test.sv