../../common/tb/prover_interpolate_cubic_test.sv