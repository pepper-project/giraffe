../../common/rtl/verifier_adder_tree.sv