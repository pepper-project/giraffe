../../common/rtl/verifier_compute_beta_elem.sv