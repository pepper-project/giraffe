../../common/tb/prover_interpolate_qc_test.sv