../../common/tb/verifier_compute_wpreds_test.sv