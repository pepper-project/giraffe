../../common/rtl/prover_compute_v_sr.sv