../../common/func/func_lvlNumInputs.sv