../../common/rtl/prover_shim.sv